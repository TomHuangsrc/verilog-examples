module sub_module3 (
    input wire clk,
    input wire rst,
    output wire out
);

	// Some logic here
endmodule