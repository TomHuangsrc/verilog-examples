module sub_module2 (
    input wire clk,
    input wire rst,
    output wire out
);
    // Some logic here
endmodule