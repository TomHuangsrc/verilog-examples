`timescale 1ns/1ps
module sim_top_tb();

reg clk;
reg rst;

reg valid_desc;
reg [511:0] data_desc;

reg valid_qual;
reg [511:0] data_qual;

reg   item_start;
wire [7:0]       row;
wire [7:0]       col;
wire [15:0]      start_addr;
wire [7:0]       length;

assign          row=DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_waddr_f1p1[11:5];
assign          col=DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_waddr_f1p1[4:0];
assign          start_addr=DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_din_f1p1[23:16]*32+DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_din_f1p1[15:8];
assign          length=DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_din_f1p1[7:0];

integer       handle,tuple_file,item_file;

initial
begin
   handle    =$fopen("ram_index.txt");
   tuple_file=$fopen("tuple_file.txt");	
   item_file =$fopen("item_file.txt");	
end 
//divide tuple inform into detail
always@(negedge clk)
begin
   if(DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_wr_f1p1==1'd1)begin
        $fdisplay(handle,"row=%h,col=%h,addr=%h,length=%h",row,col,start_addr,length);
   end	
end
//item of tuple decode
always@(posedge clk) begin			  			
		if(DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_wr_f1p1==1'd1)
	   $fwrite(tuple_file,"addr=%h,din=%h\n",DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_waddr_f1p1,DUT.acc_engine_u1.item_unit.tuple_decode_inst.tuple_ram_din_f1p1);	

end
//the output of item decode
always@(posedge clk) begin			  			
		if(DUT.acc_engine_u1.item_unit.item_decode_inst.ram_index_wr_r==1'd1)
			$fwrite(item_file,"addr=%h,din=%h\n",DUT.acc_engine_u1.item_unit.item_decode_inst.ram_index_addr_r,DUT.acc_engine_u1.item_unit.item_decode_inst.ram_index_data_r);	

end	

    initial begin
    clk = 0;
		forever
		#5 clk = ~clk;
	end
	initial
		begin
		tuple_file=$fopen("tuple_file.txt");		
		end	
		
	initial begin
			rst = 1;
            #500;            			
		    rst = 0;	
	end

    initial begin
			valid_desc   = 1'b0;
			data_desc  = 512'b0;	
            valid_qual   = 1'b0;
			data_qual  = 512'b0;
           	item_start =1'b0;		
		
	  #2000; // update key 1st
	  @(negedge clk);
	    #10;
	         valid_desc   = 1;
		     data_desc= 512'h00000000000000000000000000000000000079656b726564726f5f6c0000401600007f4013d23820000000000000000200000000ffffffff0000401800000010;
        #10; data_desc= 512'h01697001ffffffff000000000000000000010004ffffffff00000017000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h000000000000000000000000000000000000000000000000000000000000000000000079656b747261705f6c0000401600000000000000000000000100000000;
        #10; data_desc= 512'h0000000000000000000000010000000001697001ffffffffffffffff0000000000020004ffffffff000000170000000000000000000000000000000000000000;
        #10; data_desc= 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000079656b707075735f6c00004016;
        #10; data_desc= 512'h7265626d756e656e696c5f6c000040160000000000000000000000010000000001697001ffffffffffffffff0000000000030004ffffffff0000001700000000;
        #10; data_desc= 512'h00040004ffffffff0000001700000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h000000000000000000000000000000000000797469746e6175715f6c000040160000000000000000000000010000000001697001ffffffffffffffff00000000;
        #10; data_desc= 512'h01647001ffffffffffffffff0000000000050008ffffffff000002bd000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h000000000000000000000000000000000000000000000000000000000065636972706465646e657478655f6c0000401600000000000000000000000100000000;
        #10; data_desc= 512'h0000000000000000000000010000000001647001ffffffffffffffff0000000000060008ffffffff000002bd0000000000000000000000000000000000000000;
        #10; data_desc= 512'h0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000746e756f637369645f6c00004016;
        #10; data_desc= 512'h000000000000007861745f6c000040160000000000000000000000010000000001647001ffffffffffffffff0000000000070008ffffffff000002bd00000000;
        #10; data_desc= 512'h00080008ffffffff000002bd00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h0000000000000000000000000000000067616c666e72757465725f6c000040160000000000000000000000010000000001647001ffffffffffffffff00000000;
        #10; data_desc= 512'h0169700000000005ffffffff000000000009ffffffffffff00000412000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h0000000000000000000000000000000000000000000000000000000000000000737574617473656e696c5f6c0000401600000064000000000000000100000000;
        #10; data_desc= 512'h000000640000000000000001000000000169700000000005ffffffff00000000000affffffffffff000004120000000000000000000000000000000000000000;
        #10; data_desc= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000065746164706968735f6c00004016;
        #10; data_desc= 512'h6574616474696d6d6f635f6c000040160000000000000000000000010000000001697001ffffffffffffffff00000000000b0004ffffffff0000043a00000000;
        #10; data_desc= 512'h000c0004ffffffff0000043a00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h00000000000000000000000000000065746164747069656365725f6c000040160000000000000000000000010000000001697001ffffffffffffffff00000000;
        #10; data_desc= 512'h01697001ffffffffffffffff00000000000d0004ffffffff0000043a000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h0000000000000000000000000000000000000000000000000000000000007463757274736e69706968735f6c0000401600000000000000000000000100000000;
        #10; data_desc= 512'h00000064000000000000000100000000016970000000001dffffffff00000000000effffffffffff000004120000000000000000000000000000000000000000;
        #10; data_desc= 512'h000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000065646f6d706968735f6c00004016;
        #10; data_desc= 512'h000000746e656d6d6f635f6c0000401600000064000000000000000100000000016970000000000effffffff00000000000fffffffffffff0000041200000000;
        #10; data_desc= 512'h0010ffffffffffff0000041300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h0000000000000000000000000000000000000000000000000000000000000000000000640000000000000001000000000169700000000030ffffffff00000000;   //real end
		#10; data_desc= 512'h0010ffffffffffff0000041300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_desc= 512'h0000000000000000000000000000000000000000000000000000000000000000000000640000000000000001000000000169700000000030ffffffff00000000;
        #10; valid_desc = 0; 		//memcpy_done
		     data_desc  =512'b0;
		#1000;
	    #10;
	         valid_qual   = 1;
             data_qual = 512'h71010000000a028b0000044049000000000000020100000000000000040102850000043fa999999999999a0201000000000000000601028b0000003022030102;
        #10; data_qual = 512'hde010000000a02850000000000000000000000000000000000000000000000000000143fb1eb851eb851ec0201000000000000000601028c0000000004fffff7;
        #10; data_qual = 512'h00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000587631302011100581080000000014fffff8; //read end
		#10; data_qual = 512'h0010ffffffffffff0000041300000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000;
        #10; data_qual = 512'h0000000000000000000000000000000000000000000000000000000000000000000000640000000000000001000000000169700000000030ffffffff00000000;
        #10; valid_qual  = 0; 		//memcpy_done
		     data_qual =512'b0;
			 
		#2000;
             item_start=1'b1;
		#10;
		     item_start=1'b0;
    end
sim_top DUT(
.clk(clk),
.rst(rst),

.item_start(item_start),

.rdata_reg_desc  (data_desc),
.rvalid_reg_desc (valid_desc),

.rdata_reg_qual  (data_qual),
.rvalid_reg_qual (valid_qual)
);

endmodule
